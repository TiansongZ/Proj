//second version
